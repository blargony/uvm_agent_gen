{% extends "_base.sv" %}

{% block body %}

`include "{{ agent.name }}_nominal_seq.sv"

{% endblock %}
